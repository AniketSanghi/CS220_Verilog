`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:10:28 02/06/2019 
// Design Name: 
// Module Name:    printstring 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module printstring(LCD_E, LCD_RS, LCD_W, data);

output LCD_E, LCD_RS, LCD_W;
output [3:0] data;


endmodule
